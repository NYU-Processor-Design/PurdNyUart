module Uart;

endmodule
